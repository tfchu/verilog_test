`include "test.sv"

module top
    initial begin
        run_test("feature_test");
    end
endmodule
`define NUM_BITS 4


program automatic test;
    initial begin
        $display(`NUM_BITS);

    end
endprogram 
/**

// no monitor and scoreboard
[ DRIVER ] ----- Reset Started -----
[ DRIVER ] ----- Reset Ended   -----
-------------------------
- [ Generator ] 
-------------------------
- a = 13, b = 2
- c = 0
-------------------------
-------------------------
- [ Generator ] 
-------------------------
- a = 6, b = 4
- c = 0
-------------------------
-------------------------
- [ Generator ] 
-------------------------
- a = 15, b = 11
- c = 0
-------------------------
-------------------------
- [ Generator ] 
-------------------------
- a = 15, b = 5
- c = 0
-------------------------
-------------------------
- [ Driver ] 
-------------------------
- a = 13, b = 2
- c = 15
-------------------------
-------------------------
- [ Driver ] 
-------------------------
- a = 6, b = 4
- c = 10
-------------------------
-------------------------
- [ Driver ] 
-------------------------
- a = 15, b = 11
- c = 26
-------------------------
-------------------------
- [ Driver ] 
-------------------------
- a = 15, b = 5
- c = 20
-------------------------

// with monitor and scoreboard (use environment_new.sv)
[ DRIVER ] ----- Reset Started -----
[ DRIVER ] ----- Reset Ended   -----
-------------------------
- [ Generator ] 
-------------------------
- a = 13, b = 2
- c = 0
-------------------------
-------------------------
- [ Generator ] 
-------------------------
- a = 6, b = 4
- c = 0
-------------------------
-------------------------
- [ Generator ] 
-------------------------
- a = 15, b = 11
- c = 0
-------------------------
-------------------------
- [ Generator ] 
-------------------------
- a = 15, b = 5
- c = 0
-------------------------
-------------------------
- [ Driver ] 
-------------------------
- a = 13, b = 2
- c = 15
-------------------------
-------------------------
- [ Monitor ] 
-------------------------
- a = 13, b = 2
- c = 15
-------------------------
Result is as Expected
-------------------------
- [ Scoreboard ] 
-------------------------
- a = 13, b = 2
- c = 15
-------------------------
-------------------------
- [ Driver ] 
-------------------------
- a = 6, b = 4
- c = 10
-------------------------
-------------------------
- [ Monitor ] 
-------------------------
- a = 6, b = 4
- c = 10
-------------------------
Result is as Expected
-------------------------
- [ Scoreboard ] 
-------------------------
- a = 6, b = 4
- c = 10
-------------------------
-------------------------
- [ Driver ] 
-------------------------
- a = 15, b = 11
- c = 26
-------------------------
-------------------------
- [ Monitor ] 
-------------------------
- a = 15, b = 11
- c = 26
-------------------------
Result is as Expected
-------------------------
- [ Scoreboard ] 
-------------------------
- a = 15, b = 11
- c = 26
-------------------------
-------------------------
- [ Driver ] 
-------------------------
- a = 15, b = 5
- c = 20
-------------------------
-------------------------
- [ Monitor ] 
-------------------------
- a = 15, b = 5
- c = 20
-------------------------
Result is as Expected
-------------------------
- [ Scoreboard ] 
-------------------------
- a = 15, b = 5
- c = 20
-------------------------

*/

`include "interface.sv"
`include "random_test.sv"
 
module tbench_top;
   
    //clock and reset signal declaration
    bit clk;
    bit reset;
    
    //clock generation
    always #5 clk = ~clk;
    
    //reset Generation
    initial begin
        reset = 1;
        #5 reset =0;
    end
    
    //creatinng instance of interface, in order to connect DUT and testcase
    intf i_intf(clk,reset);
    
    //Testcase instance, interface handle is passed to test as an argument
    test t1(i_intf);
    
    //DUT instance, interface signals are connected to the DUT ports
    adder DUT (
        .clk(i_intf.clk),
        .reset(i_intf.reset),
        .a(i_intf.a),
        .b(i_intf.b),
        .valid(i_intf.valid),
        .c(i_intf.c)
    );
    
    //enabling the wave dump
    initial begin
        $dumpfile("dump.vcd"); $dumpvars;
    end

endmodule

/**
https://www.chipverify.com/systemverilog/systemverilog-memory-partition-constraint-example
Variable memory partitions

*/
/**
https://www.chipverify.com/systemverilog/systemverilog-memory-partition-constraint-example
Equal partitions of memory

*/
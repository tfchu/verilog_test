module not_gate(a, q);
    input  a;
    output q;

    assign q = ~a;
endmodule